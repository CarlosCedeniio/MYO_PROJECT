-- SISTEMA.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SISTEMA is
	port (
		clk_clk                        : in    std_logic                     := '0';             --                        clk.clk
		reset_reset_n                  : in    std_logic                     := '0';             --                      reset.reset_n
		sdram_addr                     : out   std_logic_vector(12 downto 0);                    --                      sdram.addr
		sdram_ba                       : out   std_logic_vector(1 downto 0);                     --                           .ba
		sdram_cas_n                    : out   std_logic;                                        --                           .cas_n
		sdram_cke                      : out   std_logic;                                        --                           .cke
		sdram_cs_n                     : out   std_logic;                                        --                           .cs_n
		sdram_dq                       : inout std_logic_vector(15 downto 0) := (others => '0'); --                           .dq
		sdram_dqm                      : out   std_logic_vector(1 downto 0);                     --                           .dqm
		sdram_ras_n                    : out   std_logic;                                        --                           .ras_n
		sdram_we_n                     : out   std_logic;                                        --                           .we_n
		sdram_clk_1_clk                : out   std_logic;                                        --                sdram_clk_1.clk
		uart_0_external_connection_rxd : in    std_logic                     := '0';             -- uart_0_external_connection.rxd
		uart_0_external_connection_txd : out   std_logic                                         --                           .txd
	);
end entity SISTEMA;

architecture rtl of SISTEMA is
	component SISTEMA_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component SISTEMA_CPU;

	component SISTEMA_JTAG is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component SISTEMA_JTAG;

	component SISTEMA_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component SISTEMA_SDRAM;

	component SISTEMA_SYS_ID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component SISTEMA_SYS_ID;

	component SISTEMA_TIMER is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component SISTEMA_TIMER;

	component SISTEMA_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component SISTEMA_pll;

	component SISTEMA_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component SISTEMA_uart_0;

	component SISTEMA_mm_interconnect_0 is
		port (
			CLOCK_clk_clk                         : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                  : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_write                 : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read           : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write             : out std_logic;                                        -- write
			CPU_debug_mem_slave_read              : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			JTAG_avalon_jtag_slave_address        : out std_logic_vector(0 downto 0);                     -- address
			JTAG_avalon_jtag_slave_write          : out std_logic;                                        -- write
			JTAG_avalon_jtag_slave_read           : out std_logic;                                        -- read
			JTAG_avalon_jtag_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_avalon_jtag_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_avalon_jtag_slave_waitrequest    : in  std_logic                     := 'X';             -- waitrequest
			JTAG_avalon_jtag_slave_chipselect     : out std_logic;                                        -- chipselect
			SDRAM_s1_address                      : out std_logic_vector(24 downto 0);                    -- address
			SDRAM_s1_write                        : out std_logic;                                        -- write
			SDRAM_s1_read                         : out std_logic;                                        -- read
			SDRAM_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                   : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                   : out std_logic;                                        -- chipselect
			SYS_ID_control_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			SYS_ID_control_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			TIMER_s1_write                        : out std_logic;                                        -- write
			TIMER_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TIMER_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			TIMER_s1_chipselect                   : out std_logic;                                        -- chipselect
			uart_0_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                       : out std_logic;                                        -- write
			uart_0_s1_read                        : out std_logic;                                        -- read
			uart_0_s1_readdata                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                   : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer               : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                  : out std_logic                                         -- chipselect
		);
	end component SISTEMA_mm_interconnect_0;

	component SISTEMA_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component SISTEMA_irq_mapper;

	component sistema_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sistema_rst_controller;

	component sistema_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component sistema_rst_controller_001;

	signal cpu_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                              : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                  : std_logic_vector(27 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                     : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_write                                    : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                           : std_logic_vector(27 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                              : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	signal mm_interconnect_0_sys_id_control_slave_readdata          : std_logic_vector(31 downto 0); -- SYS_ID:readdata -> mm_interconnect_0:SYS_ID_control_slave_readdata
	signal mm_interconnect_0_sys_id_control_slave_address           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SYS_ID_control_slave_address -> SYS_ID:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest        : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	signal mm_interconnect_0_timer_s1_readdata                      : std_logic_vector(15 downto 0); -- TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	signal mm_interconnect_0_timer_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TIMER_s1_address -> TIMER:address
	signal mm_interconnect_0_timer_s1_write                         : std_logic;                     -- mm_interconnect_0:TIMER_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                      : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                   : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                       : std_logic_vector(24 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_read                          : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                 : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                         : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_0_uart_0_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_0_uart_0_s1_readdata                     : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	signal mm_interconnect_0_uart_0_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_0_uart_0_s1_read                         : std_logic;                     -- mm_interconnect_0:uart_0_s1_read -> mm_interconnect_0_uart_0_s1_read:in
	signal mm_interconnect_0_uart_0_s1_begintransfer                : std_logic;                     -- mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_0_uart_0_s1_write                        : std_logic;                     -- mm_interconnect_0:uart_0_s1_write -> mm_interconnect_0_uart_0_s1_write:in
	signal mm_interconnect_0_uart_0_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	signal irq_mapper_receiver0_irq                                 : std_logic;                     -- TIMER:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                 : std_logic;                     -- JTAG:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                 : std_logic;                     -- uart_0:irq -> irq_mapper:receiver2_irq
	signal cpu_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                       : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                            : std_logic;                     -- CPU:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                       : std_logic;                     -- rst_controller_001:reset_out -> pll:rst
	signal reset_reset_n_ports_inv                                  : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> JTAG:av_read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> JTAG:av_write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> TIMER:write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv          : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal mm_interconnect_0_uart_0_s1_read_ports_inv               : std_logic;                     -- mm_interconnect_0_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_0_uart_0_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_uart_0_s1_write:inv -> uart_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, JTAG:rst_n, SDRAM:reset_n, SYS_ID:reset_n, TIMER:reset_n, uart_0:reset_n]

begin

	cpu : component SISTEMA_CPU
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	jtag : component SISTEMA_JTAG
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                  --               irq.irq
		);

	sdram : component SISTEMA_SDRAM
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	sys_id : component SISTEMA_SYS_ID
		port map (
			clock    => clk_clk,                                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_sys_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sys_id_control_slave_address(0)  --              .address
		);

	timer : component SISTEMA_TIMER
		port map (
			clk        => clk_clk,                                    --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                    --   irq.irq
		);

	pll : component SISTEMA_pll
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_001_reset_out_reset, --   reset.reset
			outclk_0 => sdram_clk_1_clk,                    -- outclk0.clk
			outclk_1 => open,                               -- outclk1.clk
			locked   => open                                -- (terminated)
		);

	uart_0 : component SISTEMA_uart_0
		port map (
			clk           => clk_clk,                                     --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_0_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_uart_0_s1_readdata,        --                    .readdata
			rxd           => uart_0_external_connection_rxd,              -- external_connection.export
			txd           => uart_0_external_connection_txd,              --                    .export
			irq           => irq_mapper_receiver2_irq                     --                 irq.irq
		);

	mm_interconnect_0 : component SISTEMA_mm_interconnect_0
		port map (
			CLOCK_clk_clk                         => clk_clk,                                              --                       CLOCK_clk.clk
			CPU_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                       -- CPU_reset_reset_bridge_in_reset.reset
			CPU_data_master_address               => cpu_data_master_address,                              --                 CPU_data_master.address
			CPU_data_master_waitrequest           => cpu_data_master_waitrequest,                          --                                .waitrequest
			CPU_data_master_byteenable            => cpu_data_master_byteenable,                           --                                .byteenable
			CPU_data_master_read                  => cpu_data_master_read,                                 --                                .read
			CPU_data_master_readdata              => cpu_data_master_readdata,                             --                                .readdata
			CPU_data_master_write                 => cpu_data_master_write,                                --                                .write
			CPU_data_master_writedata             => cpu_data_master_writedata,                            --                                .writedata
			CPU_data_master_debugaccess           => cpu_data_master_debugaccess,                          --                                .debugaccess
			CPU_instruction_master_address        => cpu_instruction_master_address,                       --          CPU_instruction_master.address
			CPU_instruction_master_waitrequest    => cpu_instruction_master_waitrequest,                   --                                .waitrequest
			CPU_instruction_master_read           => cpu_instruction_master_read,                          --                                .read
			CPU_instruction_master_readdata       => cpu_instruction_master_readdata,                      --                                .readdata
			CPU_debug_mem_slave_address           => mm_interconnect_0_cpu_debug_mem_slave_address,        --             CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write             => mm_interconnect_0_cpu_debug_mem_slave_write,          --                                .write
			CPU_debug_mem_slave_read              => mm_interconnect_0_cpu_debug_mem_slave_read,           --                                .read
			CPU_debug_mem_slave_readdata          => mm_interconnect_0_cpu_debug_mem_slave_readdata,       --                                .readdata
			CPU_debug_mem_slave_writedata         => mm_interconnect_0_cpu_debug_mem_slave_writedata,      --                                .writedata
			CPU_debug_mem_slave_byteenable        => mm_interconnect_0_cpu_debug_mem_slave_byteenable,     --                                .byteenable
			CPU_debug_mem_slave_waitrequest       => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,    --                                .waitrequest
			CPU_debug_mem_slave_debugaccess       => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,    --                                .debugaccess
			JTAG_avalon_jtag_slave_address        => mm_interconnect_0_jtag_avalon_jtag_slave_address,     --          JTAG_avalon_jtag_slave.address
			JTAG_avalon_jtag_slave_write          => mm_interconnect_0_jtag_avalon_jtag_slave_write,       --                                .write
			JTAG_avalon_jtag_slave_read           => mm_interconnect_0_jtag_avalon_jtag_slave_read,        --                                .read
			JTAG_avalon_jtag_slave_readdata       => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,    --                                .readdata
			JTAG_avalon_jtag_slave_writedata      => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,   --                                .writedata
			JTAG_avalon_jtag_slave_waitrequest    => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest, --                                .waitrequest
			JTAG_avalon_jtag_slave_chipselect     => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,  --                                .chipselect
			SDRAM_s1_address                      => mm_interconnect_0_sdram_s1_address,                   --                        SDRAM_s1.address
			SDRAM_s1_write                        => mm_interconnect_0_sdram_s1_write,                     --                                .write
			SDRAM_s1_read                         => mm_interconnect_0_sdram_s1_read,                      --                                .read
			SDRAM_s1_readdata                     => mm_interconnect_0_sdram_s1_readdata,                  --                                .readdata
			SDRAM_s1_writedata                    => mm_interconnect_0_sdram_s1_writedata,                 --                                .writedata
			SDRAM_s1_byteenable                   => mm_interconnect_0_sdram_s1_byteenable,                --                                .byteenable
			SDRAM_s1_readdatavalid                => mm_interconnect_0_sdram_s1_readdatavalid,             --                                .readdatavalid
			SDRAM_s1_waitrequest                  => mm_interconnect_0_sdram_s1_waitrequest,               --                                .waitrequest
			SDRAM_s1_chipselect                   => mm_interconnect_0_sdram_s1_chipselect,                --                                .chipselect
			SYS_ID_control_slave_address          => mm_interconnect_0_sys_id_control_slave_address,       --            SYS_ID_control_slave.address
			SYS_ID_control_slave_readdata         => mm_interconnect_0_sys_id_control_slave_readdata,      --                                .readdata
			TIMER_s1_address                      => mm_interconnect_0_timer_s1_address,                   --                        TIMER_s1.address
			TIMER_s1_write                        => mm_interconnect_0_timer_s1_write,                     --                                .write
			TIMER_s1_readdata                     => mm_interconnect_0_timer_s1_readdata,                  --                                .readdata
			TIMER_s1_writedata                    => mm_interconnect_0_timer_s1_writedata,                 --                                .writedata
			TIMER_s1_chipselect                   => mm_interconnect_0_timer_s1_chipselect,                --                                .chipselect
			uart_0_s1_address                     => mm_interconnect_0_uart_0_s1_address,                  --                       uart_0_s1.address
			uart_0_s1_write                       => mm_interconnect_0_uart_0_s1_write,                    --                                .write
			uart_0_s1_read                        => mm_interconnect_0_uart_0_s1_read,                     --                                .read
			uart_0_s1_readdata                    => mm_interconnect_0_uart_0_s1_readdata,                 --                                .readdata
			uart_0_s1_writedata                   => mm_interconnect_0_uart_0_s1_writedata,                --                                .writedata
			uart_0_s1_begintransfer               => mm_interconnect_0_uart_0_s1_begintransfer,            --                                .begintransfer
			uart_0_s1_chipselect                  => mm_interconnect_0_uart_0_s1_chipselect                --                                .chipselect
		);

	irq_mapper : component SISTEMA_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component sistema_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component sistema_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_uart_0_s1_read_ports_inv <= not mm_interconnect_0_uart_0_s1_read;

	mm_interconnect_0_uart_0_s1_write_ports_inv <= not mm_interconnect_0_uart_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of SISTEMA
